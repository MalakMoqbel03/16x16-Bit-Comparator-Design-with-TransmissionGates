*** SPICE deck for cell Inv_sim{lay} from library Inverter
*** Created on Fri Apr 05, 2024 15:42:03
*** Last revised on Fri Apr 05, 2024 15:44:56
*** Written on Fri Apr 26, 2024 22:58:13 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Inverter__Inv FROM CELL Inverter:Inv{lay}
.SUBCKT Inverter__Inv A gnd vdd Y
Mnmos@0 gnd A Y gnd NMOS L=0.4U W=2U AS=3P AD=8P PS=7U PD=19U
Mpmos@0 vdd A Y vdd PMOS L=0.4U W=2U AS=3P AD=9P PS=7U PD=19.4U
.ENDS Inverter__Inv

*** TOP LEVEL CELL: Inverter:Inv_sim{lay}
XInv@0 A gnd vdd Y Inverter__Inv

* Spice Code nodes in cell cell 'Inverter:Inv_sim{lay}'
vdd vdd 0 DC 5
Vin A 0 pwl 10n 0 20n 5 50n 5 60n 0
cload Y 0 250fF
.measure tran tf trig v(Y) val=4.5 fall=1 td=8ns trag v(Y) val=0.5 fall=1
.measure tran tr trig v(Y) val=0.5 rise=1 td=50ns trag v(Y) val=4.5 rise=1
.tran 0 0.1us
.include C:\electric\C5_models.txt
.END
