*** SPICE deck for cell NAND{lay} from library 3_Input_NAND
*** Created on Fri Apr 26, 2024 19:04:52
*** Last revised on Sat Apr 27, 2024 02:04:49
*** Written on Sat Apr 27, 2024 02:05:15 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: 3_Input_NAND:NAND{lay}
Mnmos@0 gnd X1 net@0 gnd NMOS L=0.4U W=2U AS=1P AD=10P PS=3U PD=23U
Mnmos@1 net@0 X2 net@2 gnd NMOS L=0.4U W=2U AS=0.79P AD=1P PS=3U PD=3U
Mnmos@2 net@2 X3 Y gnd NMOS L=0.4U W=2U AS=2.55P AD=0.79P PS=5.55U PD=3U
Mpmos@0 vdd X1 Y vdd PMOS L=0.4U W=2U AS=2.55P AD=4.733P PS=5.55U PD=10.733U
Mpmos@1 Y X2 vdd vdd PMOS L=0.4U W=2U AS=4.733P AD=2.55P PS=10.733U PD=5.55U
Mpmos@2 vdd X3 Y vdd PMOS L=0.4U W=2U AS=2.55P AD=4.733P PS=5.55U PD=10.733U

* Spice Code nodes in cell cell '3_Input_NAND:NAND{lay}'
vdd vdd 0 DC 5
Vx1 X1 0 pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
Vx2 X2 0 pwl 10n 0 20n 5 100n 5 110n 0
Vx3 X3 0 pwl 10n 0 20n 5 150n 5 160n 0
cload Y 0 375fF
.measure tran tf trig v(Y) val=4.5 fall=1 td=4ns trag v(Y) val=0.5 fall=1
.measure tran tr trig v(Y) val=0.5 rise=1 td=4ns trag v(Y) val=4.5 rise=1
.tran 200n
.include C:\electric\C5_models.txt 
.END
