*** SPICE deck for cell NOR{lay} from library 3_Input_NOR
*** Created on Sat Apr 27, 2024 04:18:38
*** Last revised on Sat Apr 27, 2024 06:02:14
*** Written on Sat Apr 27, 2024 06:42:39 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: 3_Input_NOR:NOR{lay}
Mnmos@0 gnd X1 Y gnd NMOS L=0.4U W=2U AS=2.4P AD=5P PS=5.4U PD=11U
Mnmos@1 Y X2 gnd gnd NMOS L=0.4U W=2U AS=5P AD=2.4P PS=11U PD=5.4U
Mnmos@2 gnd X3 Y gnd NMOS L=0.4U W=2U AS=2.4P AD=5P PS=5.4U PD=11U
Mpmos@0 vdd X1 net@0 vdd PMOS L=0.4U W=2U AS=1.2P AD=12.6P PS=3.2U PD=25.4U
Mpmos@1 net@0 X2 net@1 vdd PMOS L=0.4U W=2U AS=1P AD=1.2P PS=3U PD=3.2U
Mpmos@2 net@1 X3 Y vdd PMOS L=0.4U W=2U AS=2.4P AD=1P PS=5.4U PD=3U

* Spice Code nodes in cell cell '3_Input_NOR:NOR{lay}'
vdd vdd 0 DC 5
Vx1 X1 0 pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
Vx2 X2 0 pwl 10n 0 20n 5 100n 5 110n 0
Vx3 X3 0 pwl 10n 0 20n 5 150n 5 160n 0
cload Y 0 375fF
.measure tran tf trig v(Y) val=4.5 fall=1 td=4ns trag v(Y) val=0.5 fall=1
.measure tran tr trig v(Y) val=0.5 rise=1 td=4ns trag v(Y) val=4.5 rise=1
.tran 200n
.include C:\electric\C5_models.txt 
.END
