*** SPICE deck for cell 1bit{sch} from library 1bit
*** Created on Tue May 28, 2024 01:36:55
*** Last revised on Tue May 28, 2024 01:45:39
*** Written on Tue May 28, 2024 01:45:48 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Inverter__Inv FROM CELL Inverter:Inv{sch}
.SUBCKT Inverter__Inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=0.6U W=3U
Mpmos@0 vdd in out vdd PMOS L=0.6U W=3U
.ENDS Inverter__Inv

*** SUBCIRCUIT _3_Input_NAND__NAND FROM CELL 3_Input_NAND:NAND{sch}
.SUBCKT _3_Input_NAND__NAND X1 X2 Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y X1 net@16 gnd NMOS L=0.6U W=1.8U
Mnmos@1 net@16 X2 gnd gnd NMOS L=0.6U W=1.8U
Mpmos@1 vdd X2 Y vdd PMOS L=0.6U W=3.6U
Mpmos@2 vdd X1 Y vdd PMOS L=0.6U W=3.6U
.ENDS _3_Input_NAND__NAND

*** SUBCIRCUIT NOR2__NOR2 FROM CELL NOR2:NOR2{sch}
.SUBCKT NOR2__NOR2 X1 X2 Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 Y X1 gnd gnd NMOS L=0.6U W=1.8U
Mnmos@2 Y X2 gnd gnd NMOS L=0.6U W=1.8U
Mpmos@1 vdd X1 net@20 vdd PMOS L=0.6U W=3.6U
Mpmos@2 net@20 X2 Y vdd PMOS L=0.6U W=3.6U
.ENDS NOR2__NOR2

.global gnd vdd

*** TOP LEVEL CELL: 1bit{sch}
XInv@0 A net@5 Inverter__Inv
XInv@1 net@28 ABprime Inverter__Inv
XInv@2 net@8 AprimeB Inverter__Inv
XInv@3 B net@19 Inverter__Inv
XNAND@0 net@5 B net@28 _3_Input_NAND__NAND
XNAND@1 A net@19 net@8 _3_Input_NAND__NAND
XNOR2@2 ABprime AprimeB EQ NOR2__NOR2

* Spice Code nodes in cell cell '1bit{sch}'
vdd vdd 0 DC 5
Vx1 B 0 pwl 10n 0 20n 5 30n 5 40n 0 60n 0 
Vx2 A 0 pwl 10n 0 20n 0 30n 0 40n 5 60n 0
cload ABprime 0 375fF
cload1 AprimeB 0 375fF
cload2 EQ 0 375fF
.measure tran tf trig v(ABprime) val=4.5 fall=1 td=4ns trag v(ABprime) val=0.5 fall=1
.measure tran tr trig v(ABprime) val=0.5 rise=1 td=4ns trag v(ABprime) val=4.5 rise=1
.measure tran tf1 trig v(AprimeB) val=4.5 fall=1 td=4ns trag v(AprimeB) val=0.5 fall=1
.measure tran tr1 trig v(AprimeB) val=0.5 rise=1 td=4ns trag v(AprimeB) val=4.5 rise=1
.measure tran tf2 trig v(EQ) val=4.5 fall=1 td=4ns trag v(EQ) val=0.5 fall=1
.measure tran tr2 trig v(EQ) val=0.5 rise=1 td=4ns trag v(EQ) val=4.5 rise=1
.tran 200n
.include C:\electric\C5_models.txt
.END
