*** SPICE deck for cell Inv_sch{sch} from library Inverter
*** Created on Thu Apr 04, 2024 15:51:53
*** Last revised on Fri Apr 05, 2024 15:44:23
*** Written on Fri Apr 05, 2024 15:44:32 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Inverter__Inv FROM CELL Inv{sch}
.SUBCKT Inverter__Inv A Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y A gnd gnd NMOS L=0.4U W=2U
Mpmos@0 vdd A Y vdd PMOS L=0.4U W=2U
.ENDS Inverter__Inv

.global gnd vdd

*** TOP LEVEL CELL: Inv_sch{sch}
XInv@0 A Y Inverter__Inv

* Spice Code nodes in cell cell 'Inv_sch{sch}'
vdd vdd 0 DC 5
Vin A 0 pwl 10n 0 20n 5 50n 5 60n 0
cload Y 0 250fF
.measure tran tf trig v(Y) val=4.5 fall=1 td=8ns trag v(Y) val=0.5 fall=1
.measure tran tr trig v(Y) val=0.5 rise=1 td=50ns trag v(Y) val=4.5 rise=1
.tran 0 0.1us
.include C:\electric\C5_models.txt
.END
