*** SPICE deck for cell 2-bit_Comparator{sch} from library 2-bit_Comparator
*** Created on Thu May 30, 2024 18:18:19
*** Last revised on Sat Jun 15, 2024 15:35:53
*** Written on Sat Jun 15, 2024 15:41:01 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Inverter__Inv FROM CELL Inverter:Inv{sch}
.SUBCKT Inverter__Inv A Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y A gnd gnd NMOS L=0.4U W=2U
Mpmos@0 vdd A Y vdd PMOS L=0.4U W=2U
.ENDS Inverter__Inv

*** SUBCIRCUIT _2_Input_NAND__NAND FROM CELL 2_Input_NAND:NAND{sch}
.SUBCKT _2_Input_NAND__NAND X1 X2 Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y X1 net@16 gnd NMOS L=0.4U W=1.2U
Mnmos@1 net@16 X2 gnd gnd NMOS L=0.4U W=1.2U
Mpmos@1 vdd X2 Y vdd PMOS L=0.4U W=2.4U
Mpmos@2 vdd X1 Y vdd PMOS L=0.4U W=2.4U
.ENDS _2_Input_NAND__NAND

*** SUBCIRCUIT _2_Input_NOR__NOR FROM CELL 2_Input_NOR:NOR{sch}
.SUBCKT _2_Input_NOR__NOR X2 X3 Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y X3 Y gnd NMOS L=0.4U W=1.2U
Mnmos@1 Y X2 gnd gnd NMOS L=0.4U W=1.2U
Mpmos@1 vdd X2 net@2 vdd PMOS L=0.4U W=2.4U
Mpmos@2 net@2 X3 Y vdd PMOS L=0.4U W=2.4U
.ENDS _2_Input_NOR__NOR

*** SUBCIRCUIT _1-bit_Comparator__1-bit_Comparator FROM CELL 1-bit_Comparator:1-bit_Comparator{sch}
.SUBCKT _1-bit_Comparator__1-bit_Comparator A ABprime AprimeB B EQ
** GLOBAL gnd
** GLOBAL vdd
XInv@0 B net@1 Inverter__Inv
XInv@1 net@0 ABprime Inverter__Inv
XInv@2 net@18 AprimeB Inverter__Inv
XInv@3 A net@4 Inverter__Inv
XNAND@0 net@1 A net@0 _2_Input_NAND__NAND
XNAND@1 B net@4 net@18 _2_Input_NAND__NAND
XNOR@0 ABprime AprimeB EQ _2_Input_NOR__NOR
.ENDS _1-bit_Comparator__1-bit_Comparator

.global gnd vdd

*** TOP LEVEL CELL: 2-bit_Comparator:2-bit_Comparator{sch}
X_1-bit_Co@0 A1 net@68 net@76 B1 net@15 _1-bit_Comparator__1-bit_Comparator
X_1-bit_Co@1 A0 net@27 net@61 B0 net@12 _1-bit_Comparator__1-bit_Comparator
XInv@0 net@9 EQ Inverter__Inv
XInv@1 net@30 net@62 Inverter__Inv
XInv@2 net@69 A>B Inverter__Inv
XInv@3 net@57 B>A Inverter__Inv
XInv@4 net@50 net@72 Inverter__Inv
XNAND@0 net@15 net@12 net@9 _2_Input_NAND__NAND
XNAND@1 net@15 net@27 net@30 _2_Input_NAND__NAND
XNAND@2 net@61 net@15 net@50 _2_Input_NAND__NAND
XNOR@0 net@68 net@62 net@69 _2_Input_NOR__NOR
XNOR@1 net@72 net@76 net@57 _2_Input_NOR__NOR

* Spice Code nodes in cell cell '2-bit_Comparator:2-bit_Comparator{sch}'
vdd vdd 0 DC 5
* Input signals for 2-bit comparator
Vx1 B1 0 pwl 10n 5 50n 5 90n 0 140n 0 200n 0
Vx2 A1 0 pwl 10n 0 50n 5 90n 5 140n 0 200n 0
Vx3 B0 0 pwl 10n 0 50n 0 90n 0 140n 5 200n 5
Vx4 A0 0 pwl 10n 0 50n 5 90n 5 140n 0 200n 0
cload A>B 0 375fF
cload1 B>A 0 375fF
cload2 EQ 0 375fF
.measure tran tf trig v(A>B) val=4.5 fall=1 td=4ns trag v(A>B) val=0.5 fall=1
.measure tran tr trig v(A>B) val=0.5 rise=1 td=4ns trag v(A>B) val=4.5 rise=1
.measure tran tf1 trig v(B>A) val=4.5 fall=1 td=4ns trag v(B>A) val=0.5 fall=1
.measure tran tr1 trig v(B>A) val=0.5 rise=1 td=4ns trag v(B>A) val=4.5 rise=1
.measure tran tf2 trig v(EQ) val=4.5 fall=1 td=4ns trag v(EQ) val=0.5 fall=1
.measure tran tr2 trig v(EQ) val=0.5 rise=1 td=4ns trag v(EQ) val=4.5 rise=1
.tran 200n
.include C:\electric\C5_models.txt
.END
